`default_nettype none
//a single inverter
module tt_inv (
	input  wire a,
         output wire y);

	not (y, a);

endmodule 
